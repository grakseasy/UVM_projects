class fifo_master_sequence extends uvm_sequence#(fifo_transaction);  

  `uvm_object_utils(fifo_master_sequence)

  function new (string name = "");
    super.new(name);
  endfunction

  task body();
	       repeat(12) begin
		  `uvm_do_with(req, { req.wr_en == 1; req.rd_en == 0; })
	       end
  endtask

endclass

