class master_monitor extends uvm_monitor;
  
  `uvm_component_utils(master_monitor)
  
  virtual interf vintf;
  fifo_transaction fifo_trans;
  uvm_analysis_port #(fifo_transaction) ip;

  
  function new(string name, uvm_component parent);
    super.new(name,parent);
    fifo_trans = new();
    ip = new("ip", this);
    `uvm_info("master monitor", $sformatf("Monitor: Input"), UVM_HIGH)
  endfunction
  
 function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual interf)::get(this,"","vintf",vintf)) begin
      `uvm_error("","uvm_get_config interface failed\n");
    end
  endfunction
   
  virtual task run_phase(uvm_phase phase);
     super.run_phase(phase);
     fork
		begin
		 	`uvm_info("master monitor", $sformatf("Monitor: Input\n"), UVM_HIGH)
		 	forever begin
				fifo_trans=fifo_transaction::type_id::create("fifo_trans");
			 	@(posedge vintf.clk);
				if(vintf.wr_en && !vintf.rd_en && vintf.rst)
					begin
						fifo_trans.din = vintf.din;
						fifo_trans.wr_en = vintf.wr_en;
						fifo_trans.rd_en = vintf.rd_en;
						fifo_trans.empty = vintf.empty;
						fifo_trans.wrap_on_full = vintf.wrap_on_full;
						fifo_trans.full = vintf.full;
						ip.write(fifo_trans);
						`uvm_info("MASTER MONITOR", $sformatf("MONITOR: Input = %0h", fifo_trans.din), UVM_HIGH)
					end
				if(vintf.full)
					begin
						fifo_trans.full = vintf.full;
						ip.write(fifo_trans);	
					end
			end
		end
		begin
			//reset not needed
		end
     join
  endtask
endclass
       
       
       
