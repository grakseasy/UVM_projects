package ahb_pkg;
 import uvm_pkg::*;
`include "uvm_macros.svh"
`include "transaction.sv"
`include "master_sequence.sv"
`include "sequencer.sv"
`include "master_driver.sv"
`include "master_monitor.sv"
`include "master_agent.sv"
`include "slave_sequence.sv"
`include "slave_driver.sv"
`include "slave_monitor.sv"
`include "slave_agent.sv"
`include "ahb_coverage.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"


endpackage
