package fifo_pkg;
 import uvm_pkg::*;
`include "uvm_macros.svh"

`include "fifo_transaction.sv"
`include "fifo_master_sequence.sv"
`include "fifo_master_driver.sv"
`include "fifo_master_monitor.sv"
`include "fifo_slave_sequence.sv"
`include "fifo_slave_driver.sv"
`include "fifo_slave_monitor.sv"
`include "fifo_master_agent.sv"
`include "fifo_slave_agent.sv"
`include "fifo_cov.sv"
`include "scoreboard.sv"
`include "fifo_env.sv"
`include "fifo_test.sv"


endpackage
